.SUBCKT LM317_TI in adj out
* PEI 08/98 p62
J1 in out 4 JN
Q2 5 5 6 QPL .1
Q3 5 8 9 QNL .2
Q4 8 5 7 QPL .1
Q5 81 8 out QNL .2
Q6 out 81 10 QPL .2
Q7 12 81 13 QNL .2
*Q8 10 5 11 QPL .2
Q8 A10 5 11 QPL .2
Q9 14 12 10 QPL .2
Q10 16 5 17 QPL .2
Q11 16 14 15 QNL .2 OFF
Q12 out 20 16 QPL .2
Q13 in 19 20 QNL .2
Q14 19 5 18 QPL .2
Q15 out 21 19 QPL .2
Q16 21 22 16 QPL .2
Q17 21 out 24 QNL .2
Q18 22 22 16 QPL .2
Q19 22 out 241 QNL .2
Q20 out 25 16 QPL .2
Q21 25 26 out QNL .2
Q22A 35 35 in QPL .2
Q22B 16 35 in QPL .2
Q23 35 16 30 QNL .2
Q24A 27 40 29 QNL .2
Q24B 27 40 28 QNL .2
Q25 in 31 41 QNL 5
Q26 in 41 32 QNL 50
D1 out 4 DZ
D2 33 in DZ
D3 29 34 DZ
R1 in 6 310
R2 in 7 310
R3 in 11 190
R4 in 17 82
R5 in 18 5.6K
R6 4 8 100K
R7 8 81 130
*R8 10 12 12.4K
R8 A10 12 12.4K
R9 9 out 180
R10 13 out 4.1K
R11 14 out 5.8K
R12 15 out 72
R13 20 out 5.1K
R14 adj 24 12K
R15 24 241 2.4K
R16 16 25 6.7K
R17 16 40 12K
R18 30 41 130
R19 16 31 370
R20 26 27 13K
R21 27 40 400
R22 out 41 160
R23 33 34 18K
R24 28 29 160
R25 28 32 3
R26 32 out .1
C1 21 out 30PF
C2 21 adj 30PF
C3 25 26 5PF
CBS1 5 out 2PF
CBS2 35 out 1PF
CBS3 22 out 1PF
.MODEL JN NJF (BETA=1E-4 VTO=-7)
.MODEL DZ D(BV=6.3)
.MODEL QNL NPN (EG=1.22 BF=80 RB=100 CCS=1.5PF TF=.3NS TR=6NS
+ CJE=2PF CJC=1PF VAF=100 IS=1E-22 NF=1.2)
.MODEL QPL PNP (BF=40 RB=20 TF=.6NS TR=10NS CJE=1.5PF CJC=1PF VAF=50
+ IS=1E-22 NF=1.2)
.ENDS LM317_TI